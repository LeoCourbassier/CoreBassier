module InstructionsMemory
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=10)
(
	input [(ADDR_WIDTH-1):0] read_addr,
	input clk,
	output reg [(DATA_WIDTH-1):0] q
);

	// Declare the RAM variable
	reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];

	initial 
	begin
		$readmemb("inst.txt", ram);
		// Fibonacci
		/*ram[0] = 32'b01110100001000000000000000000000;
		ram[1] = 32'b00000100010000000000000000000001;
		ram[2] = 32'b00000000011000100000100000000000;
		ram[3] = 32'b01101100110000000000000000000000;
		ram[4] = 32'b00000100101000000000000000000011;
		ram[5] = 32'b01110100001000100000000000000000;
		ram[6] = 32'b01110100010000110000000000000000;
		ram[7] = 32'b00000000011000100000100000000000;
		ram[8] = 32'b00000100101001010000000000000001;
		ram[9] = 32'b00100100111001010011000000000000;
		ram[10] = 32'b00000101000000000000000000000001;
		ram[11] = 32'b01011100111010000000000000000101;
		ram[12] = 32'b01100100000000000000000000000000;
		ram[13] = 32'b01110000000000110000000000000000;
		ram[14] = 32'b01101000000000000000000000000000;*/

		// Fatorial
		/*ram[0] = 32'b01101100110000000000000000000000;
		ram[1] = 32'b00000100001000000000000000000001;
		ram[2] = 32'b00000100010000000000000000000001;
		ram[3] = 32'b00010000010000100000100000000000;
		ram[4] = 32'b00000100001000010000000000000001;
		ram[5] = 32'b01001000011000010011000000000000;
		ram[6] = 32'b01011100000000110000000000000011;
		ram[7] = 32'b01011000000000000000000000001010;
		ram[8] = 32'b01100100000000000000000000000000;
		ram[9] = 32'b01100100000000000000000000000000;
		ram[10] = 32'b01100100000000000000000000000000;
		ram[11] = 32'b01110000000000100000000000000000;
		ram[12] = 32'b01101000000000000000000000000000;*/

		// Input to memory
		/*ram[0] = 32'b01101100010000000000000000000000;
		ram[1] = 32'b01010100000000100000000000000000;
		ram[2] = 32'b01010000011000000000000000000000;
		ram[3] = 32'b01110000000000110000000000000000;
		ram[4] = 32'b01101000000000000000000000000000;*/
	end

	always @ (posedge clk)
	begin
		q <= ram[read_addr];
	end
endmodule
