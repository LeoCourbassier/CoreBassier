module main(
				clock, sw0, sw1, sw2, sw3, sw4, sw5, sw6, sw7, sw8, sw9, sw10, sw11, sw12, sw13, sw14, sw15, sw16, sw17, 
				key0, key1, key2, key3,
				hex0, hex1, hex2, hex3, hex4, hex5, hex6, hex7,
	/*			clock2
    , halt
    , _programCounter,
    , instructionOut,
	, aluCode,
    , targetRegister, aluSource,
    , writeRegister, memoryWrite, memoryRead, memoryToRegister, branch,
    , immediate,
    , branchSignal,
    , aluBranchSignal,
    , dataA, dataB,
    , dataToWrite,
	, aluSource1, aluSource2,
    , aluError,
    , aluOut,
    , error, overflow,
	 , jump
    , memoryOut,
    inputOut,
    makeIO*/
    );

    // Inputs
    input clock;
    input sw0, sw1, sw2, sw3, sw4, sw5, sw6, sw7, sw8, sw9, sw10, sw11, sw12, sw13, sw14, sw15, sw16, sw17;
    input key0, key1, key2, key3;

    // Temporary
    wire clock2;
    wire halt;
    wire [31:0] _programCounter;
	wire [31:0] instructionOut;
	wire [5:0] aluCode;
    wire targetRegister, aluSource;
    wire writeRegister, memoryWrite, memoryRead;
    wire [2:0] memoryToRegister;
    wire branch, jump;
    reg[31:0] immediate;
    reg branchSignal;
    wire aluBranchSignal;
    wire [31:0] dataA, dataB;
    reg [31:0] dataToWrite;
	reg [31:0] aluSource1, aluSource2;
    wire aluError;
    wire [31:0] aluOut;
    wire error, overflow;
    wire [31:0] memoryOut;
    wire [31:0] inputOut;
    wire makeIO;

    // Outputs
    output [6:0] hex0, hex1, hex2, hex3, hex4, hex5, hex6, hex7;

    // Instances
    FrequencyDivider div(.clock(clock), .clockOut(clock2));
    PC programCounter(.reset(key0), .clock(clock2), .halt(halt), .immediate(immediate), .branchSignal(branchSignal), .programCounter(_programCounter), .jump(jump));
    InstructionsMemory instructionsMemory(.read_addr(_programCounter), .clk(clock2), .q(instructionOut));
    ControlUnit controlUnit(.reset(key0), .makeIO(makeIO), .clock(clock2), .opcode(instructionOut[31:26]), .aluCode(aluCode), .targetRegister(targetRegister), .aluSource(aluSource), 
        .writeRegister(writeRegister), .memoryWrite(memoryWrite), .memoryRead(memoryRead), .memoryToRegister(memoryToRegister), .branch(branch), .halt(halt), .jump(jump));
    RegistersBank registersBank(.regC(instructionOut[25:21]), 
    .regB( instructionOut[31:26] == 6'b010111 || instructionOut[31:26] == 6'b011000 ? instructionOut[25:21] : instructionOut[20:16]), 
    .regA( instructionOut[31:26] == 6'b010111 || instructionOut[31:26] == 6'b011000 ? instructionOut[20:16] : instructionOut[15:11]), 
    .writeFlag(writeRegister), .clock(clock2), .dataA(dataA), .dataB(dataB), .dataWrite(dataToWrite));
    ALU alu(.dataA(aluSource1), .dataB(aluSource2), .opCode(instructionOut[31:26]), .branchSignal(aluBranchSignal), .overflow(overflow), .error(error), .dataC(aluOut), .clock(clock2));
    DataMemory dataMemory(.data(dataB), .read_addr(aluOut), .write_addr(aluOut), .we(memoryWrite), .clk(clock), .q(memoryOut));
    IO io(.makeIO(makeIO), .reset(key0), .opcode(instructionOut[31:26]), .address(instructionOut[4:0]), .sw0(sw0), .sw1(sw1), .sw2(sw2),
     .sw3(sw3), .sw4(sw4), .sw5(sw5), .sw6(sw6), .sw7(sw7), .sw8(sw8), .sw9(sw9),
      .sw10(sw10), .sw11(sw11), .sw12(sw12), .sw13(sw13), .sw14(sw14), .sw15(sw15), .sw16(sw16),
       .sw17(sw17), .key1(key1), .key2(key2), .outL(inputOut), .hex0(hex0), 
        .hex1(hex1),  .hex2(hex2),  .hex3(hex3),  .hex4(hex4),  .hex5(hex5),  .hex6(hex6),
         .hex7(hex7), .data(dataB));
	 
    always @ ( instructionOut or aluSource or branch or aluBranchSignal or memoryToRegister )
    begin
		immediate[31:0] = { {16{instructionOut[15]}}, instructionOut[15:0] };
        branchSignal = aluBranchSignal & branch;
        
        aluSource1 = dataB;

        /* Mux for ALU input */
        case (aluSource)
            1'b0: aluSource2 = dataA;
            1'b1: aluSource2 = immediate;
        endcase

        /* Mux for writing data to register */
        case (memoryToRegister)
            3'b000: dataToWrite = aluOut;
            3'b001: dataToWrite = memoryOut;
            3'b010: dataToWrite = inputOut;
        endcase
    end
endmodule